// isp1362 device controller (D13) parameters

   parameter EPNUM_UNUSED = 12;           // number of unused endpoints

   // DC command and registers - initialization
   parameter DC_WEP0OUT_CONFIG   = 8'h20; // control endpoint OUT
   parameter DC_WEP0IN_CONFIG    = 8'h21; // control endpoint IN
   parameter DC_WEP1OUT_CONFIG   = 8'h22; // bulk endpoint OUT
   parameter DC_WEP1IN_CONFIG    = 8'h23; // bulk endpoint IN
   parameter DC_WEPNUM_CONFIG    = 8'h24; // unused endpoint starting index
   parameter DC_REP0OUT_CONIFG   = 8'h30; // control endpoint OUT
   parameter DC_REP0IN_CONIFG    = 8'h31; // control endpoint IN
   parameter DC_REP1OUT_CONIFG   = 8'h30; // bulk endpoint OUT
   parameter DC_REP1IN_CONIFG    = 8'h31; // bulk endpoint IN
   parameter DC_REPNUM_CONFIG    = 8'h32; // unused endpoint starting index
   parameter DC_WDEV_ADDR        = 8'hB6; // device address
   parameter DC_RDEV_ADDR        = 8'hB7; // address
   parameter DC_WMODE            = 8'hB8; // mode
   parameter DC_RMODE            = 8'hB9; // mode
   parameter DC_WHW_CONFIG       = 8'hBA; // hardware configuration
   parameter DC_RHW_CONIFG       = 8'hBB; // hardware configuration
   parameter DC_WIRQ_EN          = 8'hC2; // interrupt enable
   parameter DC_RIRQ_EN          = 8'hC3; // intterupt enable
   parameter DC_WRST_REG         = 8'hF6; // reset all registers
   parameter DC_WEP0OUT_BUFF     = 8'h00; // control endpoint OUT (illegal)
   parameter DC_WEP0IN_BUFF      = 8'h01; // control endpoint IN
   parameter DC_WEP1OUT_BUFF     = 8'h02; // bulk endpoint OUT (illegal)
   parameter DC_WEP1IN_BUFF      = 8'h03; // bulk endpoint IN
   parameter DC_WEPNUM_BUFF      = 8'h04; // unused endpoint starting index
   parameter DC_REP0OUT_BUFF     = 8'h10; // control endpoint OUT
   parameter DC_REP0IN_BUFF      = 8'h11; // control endpoint IN (illegal)
   parameter DC_REP1OUT_BUFF     = 8'h12; // bulk endpoint OUT
   parameter DC_REP1IN_BUFF      = 8'h13; // bulk endpoint IN
   parameter DC_REPNUM_BUFF      = 8'h14; // unused endpoint starting index
   parameter DC_SEP0OUT_STALL    = 8'h40; // control endpoint OUT (illegal)
   parameter DC_SEP0IN_STALL     = 8'h41; // control endpoint IN
   parameter DC_SEP1OUT_STALL    = 8'h42; // bulk endpoint OUT
   parameter DC_SEP1IN_STALL     = 8'h43; // bulk endpoint IN
   parameter DC_SEPNUM_STALL     = 8'h44; // endpoint starting index
   parameter DC_REP0OUT_STATUS   = 8'h50; // control endpoint OUT (illegal)
   parameter DC_REP0IN_STATUS    = 8'h51; // control endpoint IN
   parameter DC_REP1OUT_STATUS   = 8'h52; // bulk endpoint OUT
   parameter DC_REP1IN_STATUS    = 8'h53; // bulk endpoint IN
   parameter DC_REPNUM_STATUS    = 8'h54; // endpoint starting index
   parameter DC_VEP0OUT_BUFF     = 8'h60; // validate control endpoint OUT (illegal)
   parameter DC_VEP0IN_BUFF      = 8'h61; // validate control endpoint IN
   parameter DC_VEP1OUT_BUFF     = 8'h62; // validate bulk endpoint OUT
   parameter DC_VEP1IN_BUFF      = 8'h63; // validate bulk endpoint IN
   parameter DC_VEPNUM_BUFF      = 8'h64; // validate endpoint starting index
   parameter DC_CEP0OUT_BUFF     = 8'h70; // clear control endpoint OUT
   parameter DC_CEP0IN_BUFF      = 8'h71; // clear control endpoint IN (illegal)
   parameter DC_CEP1OUT_BUFF     = 8'h72; // clear bulk endpoint OUT
   parameter DC_CEP1IN_BUFF      = 8'h73; // clear bulk endpoint IN
   parameter DC_CEPNUM_BUFF      = 8'h74; // clear endpoint starting index
   parameter DC_UEP0OUT_UNSTALL  = 8'h80; // unstall control endpoint OUT (illegal)
   parameter DC_UEP0IN_UNSTALL   = 8'h81; // unstall control endpoint IN
   parameter DC_UEP1OUT_UNSTALL  = 8'h82; // unstall bulk endpoint OUT
   parameter DC_UEP1IN_UNSTALL   = 8'h83; // unstall bulk endpoint IN
   parameter DC_UEPNUM_UNSTALL   = 8'h84; // unstall endpoint starting index
   parameter DC_CHKEP0OUT_STATUS = 8'hD0; // control endpoint OUT (illegal)
   parameter DC_CHKEP0IN_STATUS  = 8'hD1; // control endpoint IN
   parameter DC_CHKEP1OUT_STATUS = 8'hD2; // bulk endpoint OUT
   parameter DC_CHKEP1IN_STATUS  = 8'hD3; // bulk endpoint IN
   parameter DC_CHKEPNUM_STATUS  = 8'hD4; // endpoint starting index
   parameter DC_ACK_SETUP        = 8'hF4; // Acknowledge Set-up EP0IN/EP0OUT
   parameter DC_REP0OUT_ERROR    = 8'hA0; // control endpoint OUT
   parameter DC_REP0IN_ERROR     = 8'hA1; // control endpoint IN
   parameter DC_REP1OUT_ERROR    = 8'hA2; // bulk endpoint OUT
   parameter DC_REP1IN_ERROR     = 8'hA3; // bulk endpoint IN
   parameter DC_REPNUM_ERROR     = 8'hA4; // unused endpoint starting index
   parameter DC_DEV_UNLOCK       = 8'hB0; // Unlock device, all registers with write access
   parameter DC_WSCRATCH_REG     = 8'hB2; // Scratch register
   parameter DC_RSCRATCH_REG     = 8'hB3; // Scratch register
   parameter DC_RFRAME_NUM       = 8'hB4; // Frame Number
   parameter DC_RCHIP_ID         = 8'hB5; // Chip ID
   parameter DC_RIRQ_REG         = 8'hC0; // Interrupt register
